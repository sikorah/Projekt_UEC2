/**
 * Copyright (C) 2024  AGH University of Science and Technology
 * MTM UEC2
 * Author: Zuzanna Schab
 *
 * Description:
 * Uart top.
 */

 module uart_top(
    input wire clk,
    input wire rst,
    input wire tx_full,
    input wire [7:0] data_second_mouse_right, 
    input wire [7:0] data_second_mouse_left, 
    output logic wr_uart,
    output logic [7:0] w_data
 );

 //local variables
logic [7:0] w_data_nxt;
logic [1:0] module_counter, module_counter_nxt;
logic wr_uart_nxt;
logic tx_tick, tx_tick_nxt;

 //logic

 always_ff @(posedge clk) begin
    if(rst) begin
        w_data <= '0;
        module_counter <= '0;
        wr_uart <= '0;
        tx_tick <= 1'b1;
    end
    else begin
        w_data <= w_data_nxt;
        module_counter <= module_counter_nxt;
        wr_uart <= wr_uart_nxt;
        tx_tick <= tx_tick_nxt;
    end
 end

 /*
 * CODES FOR MODULES
 * 00 - second_mouse_right
 * 01 - second_mouse_left
 */

 always_comb begin
    if(tx_full == 1'b0) begin
        case(module_counter)
            2'b00: begin
                w_data_nxt = data_second_mouse_right; //000
            end
            2'b01: begin
                w_data_nxt = data_second_mouse_left; //011, 100, 101, 110 
            end
           
        endcase

        if(tx_tick) begin
            module_counter_nxt = module_counter + 1;
            tx_tick_nxt = 1'b0;
        end
        else begin
            module_counter_nxt = module_counter;
            tx_tick_nxt = 1'b0;
        end
        
        if(wr_uart) begin
            wr_uart_nxt = 1'b0;
        end
        else begin
            wr_uart_nxt = 1'b1;
        end
    end
    else begin
        wr_uart_nxt = 1'b0;
        tx_tick_nxt = 1'b1;
        w_data_nxt = w_data;
        module_counter_nxt = module_counter;
    end

 end
 endmodule